import tiny8_types::*;

module tiny8v1
(
    input clk,
    input mem_resp,
    input tiny8_word mem_rdata,
    output mem_read,
    output mem_write,
    output tiny8_word mem_addr,
    output tiny8_word mem_wdata
);

/* instantiate modules here */

endmodule
