import tiny8_types::*;

module datapath
(
    input clk
);



endmodule
